* File name: D:\Documents and Settings\sicard\Mes documents\software\Dsch\Dsch35\dsch35 full\examples\amplifier\OpAmpResDivider.sch
* Software version: DSCH 3.5
* Created 19/06/2009 14:45:26
*
* Voltage and current sources
*
E1 4 0 2 3 1000
V1 7 0 DC 1.0 AC 1 0 SIN(0.0 0.5 100E6 0.0 0.0)
VDD_Div2 6 0 DC 0.5 AC 1 0
*
* Passive devices
*
R1 5 2 5K
R2 2 4 10K
R3 6 3 50
RL 8 0 50
C1 8 4 1nF
C2 5 7 1nF
*
* Active devices
*
*
* Mos models in 0.12�m
* Model 3 n-channel MOS
.MODEL  TN  NMOS
+ LEVEL=3            TPG=+1
+ GAMMA=0.2          THETA=0.5          KAPPA=0.1        ETA=0.002
+ DELTA=0.0          UO=620             VMAX=100E3       VTO=0.35
+ TOX=3e-9           XJ=0.1U            LD=0.00U         NSUB=1E+18
+ NSS=0.2            NFS=7E11
+ CJ=4.091E-4        MJ=0.307           PB=1.0
+ CJSW=3.078E-10     MJSW=1.0E-2
+ CGSO=3.93E-10      CGDO=3.93E-10
* Model 3 p-channel MOS
.MODEL  TP  PMOS
+ LEVEL=3            TPG=-1
+ GAMMA=0.2          THETA=0.5          KAPPA=0.01         ETA=0.001
+ DELTA=0.0          UO=250             VMAX=500E3         VTO=-0.35
+ TOX=3E-9          XJ=0.1U             LD=0.0U             NSUB=1E+18
+ NSS=0.0            NFS=7E11
+ CJ=6.852E-4        MJ=0.429           PB=1.0
+ CJSW=5.217E-10     MJSW=0.351
+ CGSO=7.29E-10      CGDO=7.29E-10
.TRAN 10N 10U
* Dump time and volts in "OpAmpResDivider.txt"
.control
run
set nobreak
print   V(7) V(8) V(6)  > OpAmpResDivider.txt
plot   V(7) V(8) V(6) 
.endc
.OPTIONS DELMIN=0 RELTOL=1E-6
.END
